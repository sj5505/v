module compiler

enum IntType {
	i8
	i16
	int
	i64
	i128
	byte
	u16
	u32
	u64
	u128
}

enum FloatType {
	f32
	f64
}

interface Typer{}

struct ToDo{}
